package GPIO;

module mkGPIO(Empty);
endmodule

endpackage