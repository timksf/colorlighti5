package TestHelper;
    interface TestHandler;
        method Action go();
        method Bool done();
    endinterface
endpackage
